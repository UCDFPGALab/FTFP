library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity commandInterpreter is
	port( char  : in unsigned(7 downto 0);
			readback : out std_logic);
end commandInterpreter;

architecture Behavioral of commandInterpreter is

begin


end Behavioral;

